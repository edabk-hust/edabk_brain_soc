<<<<<<< HEAD
VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO neuron_core
  CLASS BLOCK ;
  FOREIGN neuron_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 2500.000 BY 3000.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 80.590 2996.000 80.870 3000.000 ;
    END
  END clk
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 2418.310 0.000 2418.590 4.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 2986.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 2986.800 ;
    END
  END vssd1
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2468.440 2500.000 2469.040 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1594.640 4.000 1595.240 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1808.840 4.000 1809.440 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 1490.950 2996.000 1491.230 3000.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 1793.630 2996.000 1793.910 3000.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1275.040 4.000 1275.640 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2148.840 2500.000 2149.440 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1723.840 2500.000 1724.440 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 336.640 2500.000 337.240 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2128.440 4.000 2129.040 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 1713.130 0.000 1713.410 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2318.490 0.000 2318.770 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 870.440 2500.000 871.040 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 1188.270 2996.000 1188.550 3000.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2342.640 4.000 2343.240 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 582.910 2996.000 583.190 3000.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2788.040 2500.000 2788.640 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 1391.130 2996.000 1391.410 3000.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 765.040 2500.000 765.640 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1489.240 4.000 1489.840 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 1107.770 0.000 1108.050 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 955.440 4.000 956.040 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 656.240 2500.000 656.840 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1693.810 2996.000 1694.090 3000.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1914.240 4.000 1914.840 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 602.230 0.000 602.510 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 2299.170 2996.000 2299.450 3000.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 2498.810 2996.000 2499.090 3000.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1996.490 2996.000 1996.770 3000.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2573.840 2500.000 2574.440 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2893.440 2500.000 2894.040 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1404.240 2500.000 1404.840 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1190.040 2500.000 1190.640 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 685.950 2996.000 686.230 3000.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 785.770 2996.000 786.050 3000.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2363.040 2500.000 2363.640 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1088.450 2996.000 1088.730 3000.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 705.270 0.000 705.550 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 885.590 2996.000 885.870 3000.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 231.240 2500.000 231.840 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1291.310 2996.000 1291.590 3000.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2023.040 4.000 2023.640 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 483.090 2996.000 483.370 3000.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 445.440 2500.000 446.040 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2682.640 2500.000 2683.240 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 2096.310 2996.000 2096.590 3000.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 2015.810 0.000 2016.090 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1007.950 0.000 1008.230 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 975.840 2500.000 976.440 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.240 4.000 1064.840 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1383.840 4.000 1384.440 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 125.840 2500.000 126.440 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 280.230 2996.000 280.510 3000.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 2115.630 0.000 2115.910 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2553.440 4.000 2554.040 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 805.090 0.000 805.370 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 20.440 2500.000 21.040 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1615.040 2500.000 1615.640 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1084.640 2500.000 1085.240 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1915.990 0.000 1916.270 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2233.840 4.000 2234.440 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1703.440 4.000 1704.040 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.840 4.000 636.440 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1295.440 2500.000 1296.040 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2043.440 2500.000 2044.040 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2218.670 0.000 2218.950 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 2254.240 2500.000 2254.840 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1310.630 0.000 1310.910 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2767.640 4.000 2768.240 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1169.640 4.000 1170.240 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1613.310 0.000 1613.590 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 180.410 2996.000 180.690 3000.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 988.630 2996.000 988.910 3000.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2662.240 4.000 2662.840 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2199.350 2996.000 2199.630 3000.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1593.990 2996.000 1594.270 3000.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1207.590 0.000 1207.870 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2398.990 2996.000 2399.270 3000.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 550.840 2500.000 551.440 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2873.040 4.000 2873.640 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1829.240 2500.000 1829.840 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 904.910 0.000 905.190 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1410.450 0.000 1410.730 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1934.640 2500.000 1935.240 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1510.270 0.000 1510.550 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 744.640 4.000 745.240 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1896.670 2996.000 1896.950 3000.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2978.440 4.000 2979.040 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 383.270 2996.000 383.550 3000.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1812.950 0.000 1813.230 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 850.040 4.000 850.640 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2448.040 4.000 2448.640 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 2496.000 1509.640 2500.000 1510.240 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2494.120 2986.645 ;
      LAYER met1 ;
        RECT 0.070 10.640 2499.110 2986.800 ;
      LAYER met2 ;
        RECT 0.100 2995.720 80.310 2996.490 ;
        RECT 81.150 2995.720 180.130 2996.490 ;
        RECT 180.970 2995.720 279.950 2996.490 ;
        RECT 280.790 2995.720 382.990 2996.490 ;
        RECT 383.830 2995.720 482.810 2996.490 ;
        RECT 483.650 2995.720 582.630 2996.490 ;
        RECT 583.470 2995.720 685.670 2996.490 ;
        RECT 686.510 2995.720 785.490 2996.490 ;
        RECT 786.330 2995.720 885.310 2996.490 ;
        RECT 886.150 2995.720 988.350 2996.490 ;
        RECT 989.190 2995.720 1088.170 2996.490 ;
        RECT 1089.010 2995.720 1187.990 2996.490 ;
        RECT 1188.830 2995.720 1291.030 2996.490 ;
        RECT 1291.870 2995.720 1390.850 2996.490 ;
        RECT 1391.690 2995.720 1490.670 2996.490 ;
        RECT 1491.510 2995.720 1593.710 2996.490 ;
        RECT 1594.550 2995.720 1693.530 2996.490 ;
        RECT 1694.370 2995.720 1793.350 2996.490 ;
        RECT 1794.190 2995.720 1896.390 2996.490 ;
        RECT 1897.230 2995.720 1996.210 2996.490 ;
        RECT 1997.050 2995.720 2096.030 2996.490 ;
        RECT 2096.870 2995.720 2199.070 2996.490 ;
        RECT 2199.910 2995.720 2298.890 2996.490 ;
        RECT 2299.730 2995.720 2398.710 2996.490 ;
        RECT 2399.550 2995.720 2498.530 2996.490 ;
        RECT 0.100 4.280 2499.080 2995.720 ;
        RECT 0.650 3.670 99.630 4.280 ;
        RECT 100.470 3.670 199.450 4.280 ;
        RECT 200.290 3.670 299.270 4.280 ;
        RECT 300.110 3.670 402.310 4.280 ;
        RECT 403.150 3.670 502.130 4.280 ;
        RECT 502.970 3.670 601.950 4.280 ;
        RECT 602.790 3.670 704.990 4.280 ;
        RECT 705.830 3.670 804.810 4.280 ;
        RECT 805.650 3.670 904.630 4.280 ;
        RECT 905.470 3.670 1007.670 4.280 ;
        RECT 1008.510 3.670 1107.490 4.280 ;
        RECT 1108.330 3.670 1207.310 4.280 ;
        RECT 1208.150 3.670 1310.350 4.280 ;
        RECT 1311.190 3.670 1410.170 4.280 ;
        RECT 1411.010 3.670 1509.990 4.280 ;
        RECT 1510.830 3.670 1613.030 4.280 ;
        RECT 1613.870 3.670 1712.850 4.280 ;
        RECT 1713.690 3.670 1812.670 4.280 ;
        RECT 1813.510 3.670 1915.710 4.280 ;
        RECT 1916.550 3.670 2015.530 4.280 ;
        RECT 2016.370 3.670 2115.350 4.280 ;
        RECT 2116.190 3.670 2218.390 4.280 ;
        RECT 2219.230 3.670 2318.210 4.280 ;
        RECT 2319.050 3.670 2418.030 4.280 ;
        RECT 2418.870 3.670 2499.080 4.280 ;
      LAYER met3 ;
        RECT 3.990 2979.440 2496.000 2986.725 ;
        RECT 4.400 2978.040 2496.000 2979.440 ;
        RECT 3.990 2894.440 2496.000 2978.040 ;
        RECT 3.990 2893.040 2495.600 2894.440 ;
        RECT 3.990 2874.040 2496.000 2893.040 ;
        RECT 4.400 2872.640 2496.000 2874.040 ;
        RECT 3.990 2789.040 2496.000 2872.640 ;
        RECT 3.990 2787.640 2495.600 2789.040 ;
        RECT 3.990 2768.640 2496.000 2787.640 ;
        RECT 4.400 2767.240 2496.000 2768.640 ;
        RECT 3.990 2683.640 2496.000 2767.240 ;
        RECT 3.990 2682.240 2495.600 2683.640 ;
        RECT 3.990 2663.240 2496.000 2682.240 ;
        RECT 4.400 2661.840 2496.000 2663.240 ;
        RECT 3.990 2574.840 2496.000 2661.840 ;
        RECT 3.990 2573.440 2495.600 2574.840 ;
        RECT 3.990 2554.440 2496.000 2573.440 ;
        RECT 4.400 2553.040 2496.000 2554.440 ;
        RECT 3.990 2469.440 2496.000 2553.040 ;
        RECT 3.990 2468.040 2495.600 2469.440 ;
        RECT 3.990 2449.040 2496.000 2468.040 ;
        RECT 4.400 2447.640 2496.000 2449.040 ;
        RECT 3.990 2364.040 2496.000 2447.640 ;
        RECT 3.990 2362.640 2495.600 2364.040 ;
        RECT 3.990 2343.640 2496.000 2362.640 ;
        RECT 4.400 2342.240 2496.000 2343.640 ;
        RECT 3.990 2255.240 2496.000 2342.240 ;
        RECT 3.990 2253.840 2495.600 2255.240 ;
        RECT 3.990 2234.840 2496.000 2253.840 ;
        RECT 4.400 2233.440 2496.000 2234.840 ;
        RECT 3.990 2149.840 2496.000 2233.440 ;
        RECT 3.990 2148.440 2495.600 2149.840 ;
        RECT 3.990 2129.440 2496.000 2148.440 ;
        RECT 4.400 2128.040 2496.000 2129.440 ;
        RECT 3.990 2044.440 2496.000 2128.040 ;
        RECT 3.990 2043.040 2495.600 2044.440 ;
        RECT 3.990 2024.040 2496.000 2043.040 ;
        RECT 4.400 2022.640 2496.000 2024.040 ;
        RECT 3.990 1935.640 2496.000 2022.640 ;
        RECT 3.990 1934.240 2495.600 1935.640 ;
        RECT 3.990 1915.240 2496.000 1934.240 ;
        RECT 4.400 1913.840 2496.000 1915.240 ;
        RECT 3.990 1830.240 2496.000 1913.840 ;
        RECT 3.990 1828.840 2495.600 1830.240 ;
        RECT 3.990 1809.840 2496.000 1828.840 ;
        RECT 4.400 1808.440 2496.000 1809.840 ;
        RECT 3.990 1724.840 2496.000 1808.440 ;
        RECT 3.990 1723.440 2495.600 1724.840 ;
        RECT 3.990 1704.440 2496.000 1723.440 ;
        RECT 4.400 1703.040 2496.000 1704.440 ;
        RECT 3.990 1616.040 2496.000 1703.040 ;
        RECT 3.990 1614.640 2495.600 1616.040 ;
        RECT 3.990 1595.640 2496.000 1614.640 ;
        RECT 4.400 1594.240 2496.000 1595.640 ;
        RECT 3.990 1510.640 2496.000 1594.240 ;
        RECT 3.990 1509.240 2495.600 1510.640 ;
        RECT 3.990 1490.240 2496.000 1509.240 ;
        RECT 4.400 1488.840 2496.000 1490.240 ;
        RECT 3.990 1405.240 2496.000 1488.840 ;
        RECT 3.990 1403.840 2495.600 1405.240 ;
        RECT 3.990 1384.840 2496.000 1403.840 ;
        RECT 4.400 1383.440 2496.000 1384.840 ;
        RECT 3.990 1296.440 2496.000 1383.440 ;
        RECT 3.990 1295.040 2495.600 1296.440 ;
        RECT 3.990 1276.040 2496.000 1295.040 ;
        RECT 4.400 1274.640 2496.000 1276.040 ;
        RECT 3.990 1191.040 2496.000 1274.640 ;
        RECT 3.990 1189.640 2495.600 1191.040 ;
        RECT 3.990 1170.640 2496.000 1189.640 ;
        RECT 4.400 1169.240 2496.000 1170.640 ;
        RECT 3.990 1085.640 2496.000 1169.240 ;
        RECT 3.990 1084.240 2495.600 1085.640 ;
        RECT 3.990 1065.240 2496.000 1084.240 ;
        RECT 4.400 1063.840 2496.000 1065.240 ;
        RECT 3.990 976.840 2496.000 1063.840 ;
        RECT 3.990 975.440 2495.600 976.840 ;
        RECT 3.990 956.440 2496.000 975.440 ;
        RECT 4.400 955.040 2496.000 956.440 ;
        RECT 3.990 871.440 2496.000 955.040 ;
        RECT 3.990 870.040 2495.600 871.440 ;
        RECT 3.990 851.040 2496.000 870.040 ;
        RECT 4.400 849.640 2496.000 851.040 ;
        RECT 3.990 766.040 2496.000 849.640 ;
        RECT 3.990 764.640 2495.600 766.040 ;
        RECT 3.990 745.640 2496.000 764.640 ;
        RECT 4.400 744.240 2496.000 745.640 ;
        RECT 3.990 657.240 2496.000 744.240 ;
        RECT 3.990 655.840 2495.600 657.240 ;
        RECT 3.990 636.840 2496.000 655.840 ;
        RECT 4.400 635.440 2496.000 636.840 ;
        RECT 3.990 551.840 2496.000 635.440 ;
        RECT 3.990 550.440 2495.600 551.840 ;
        RECT 3.990 531.440 2496.000 550.440 ;
        RECT 4.400 530.040 2496.000 531.440 ;
        RECT 3.990 446.440 2496.000 530.040 ;
        RECT 3.990 445.040 2495.600 446.440 ;
        RECT 3.990 426.040 2496.000 445.040 ;
        RECT 4.400 424.640 2496.000 426.040 ;
        RECT 3.990 337.640 2496.000 424.640 ;
        RECT 3.990 336.240 2495.600 337.640 ;
        RECT 3.990 317.240 2496.000 336.240 ;
        RECT 4.400 315.840 2496.000 317.240 ;
        RECT 3.990 232.240 2496.000 315.840 ;
        RECT 3.990 230.840 2495.600 232.240 ;
        RECT 3.990 211.840 2496.000 230.840 ;
        RECT 4.400 210.440 2496.000 211.840 ;
        RECT 3.990 126.840 2496.000 210.440 ;
        RECT 3.990 125.440 2495.600 126.840 ;
        RECT 3.990 106.440 2496.000 125.440 ;
        RECT 4.400 105.040 2496.000 106.440 ;
        RECT 3.990 21.440 2496.000 105.040 ;
        RECT 3.990 20.040 2495.600 21.440 ;
        RECT 3.990 10.715 2496.000 20.040 ;
      LAYER met4 ;
        RECT 581.735 11.735 635.040 2985.705 ;
        RECT 637.440 11.735 711.840 2985.705 ;
        RECT 714.240 11.735 788.640 2985.705 ;
        RECT 791.040 11.735 865.440 2985.705 ;
        RECT 867.840 11.735 942.240 2985.705 ;
        RECT 944.640 11.735 1019.040 2985.705 ;
        RECT 1021.440 11.735 1095.840 2985.705 ;
        RECT 1098.240 11.735 1172.640 2985.705 ;
        RECT 1175.040 11.735 1249.440 2985.705 ;
        RECT 1251.840 11.735 1326.240 2985.705 ;
        RECT 1328.640 11.735 1403.040 2985.705 ;
        RECT 1405.440 11.735 1479.840 2985.705 ;
        RECT 1482.240 11.735 1556.640 2985.705 ;
        RECT 1559.040 11.735 1633.440 2985.705 ;
        RECT 1635.840 11.735 1710.240 2985.705 ;
        RECT 1712.640 11.735 1787.040 2985.705 ;
        RECT 1789.440 11.735 1863.840 2985.705 ;
        RECT 1866.240 11.735 1868.225 2985.705 ;
  END
END neuron_core
END LIBRARY

=======
version https://git-lfs.github.com/spec/v1
oid sha256:20796dc4843cee1414abe4e649bfd521cd092d44154975dfe6767b064de5d5af
size 32535
>>>>>>> 7fa566336ad936253585d16aa726fb716d9b4246
