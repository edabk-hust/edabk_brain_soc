version https://git-lfs.github.com/spec/v1
oid sha256:44ca5ae9246238d5a232b8f0a39fd45269beb9c97233d5fc2ba9ef1d60ae6192
size 12006
