version https://git-lfs.github.com/spec/v1
oid sha256:20796dc4843cee1414abe4e649bfd521cd092d44154975dfe6767b064de5d5af
size 32535
