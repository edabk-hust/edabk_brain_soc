magic
tech sky130A
magscale 1 2
timestamp 1699235133
<< obsli1 >>
rect 1104 2159 498824 597329
<< obsm1 >>
rect 14 2128 499822 597360
<< metal2 >>
rect 16118 599200 16174 600000
rect 36082 599200 36138 600000
rect 56046 599200 56102 600000
rect 76654 599200 76710 600000
rect 96618 599200 96674 600000
rect 116582 599200 116638 600000
rect 137190 599200 137246 600000
rect 157154 599200 157210 600000
rect 177118 599200 177174 600000
rect 197726 599200 197782 600000
rect 217690 599200 217746 600000
rect 237654 599200 237710 600000
rect 258262 599200 258318 600000
rect 278226 599200 278282 600000
rect 298190 599200 298246 600000
rect 318798 599200 318854 600000
rect 338762 599200 338818 600000
rect 358726 599200 358782 600000
rect 379334 599200 379390 600000
rect 399298 599200 399354 600000
rect 419262 599200 419318 600000
rect 439870 599200 439926 600000
rect 459834 599200 459890 600000
rect 479798 599200 479854 600000
rect 499762 599200 499818 600000
rect 18 0 74 800
rect 19982 0 20038 800
rect 39946 0 40002 800
rect 59910 0 59966 800
rect 80518 0 80574 800
rect 100482 0 100538 800
rect 120446 0 120502 800
rect 141054 0 141110 800
rect 161018 0 161074 800
rect 180982 0 181038 800
rect 201590 0 201646 800
rect 221554 0 221610 800
rect 241518 0 241574 800
rect 262126 0 262182 800
rect 282090 0 282146 800
rect 302054 0 302110 800
rect 322662 0 322718 800
rect 342626 0 342682 800
rect 362590 0 362646 800
rect 383198 0 383254 800
rect 403162 0 403218 800
rect 423126 0 423182 800
rect 443734 0 443790 800
rect 463698 0 463754 800
rect 483662 0 483718 800
<< obsm2 >>
rect 20 599144 16062 599298
rect 16230 599144 36026 599298
rect 36194 599144 55990 599298
rect 56158 599144 76598 599298
rect 76766 599144 96562 599298
rect 96730 599144 116526 599298
rect 116694 599144 137134 599298
rect 137302 599144 157098 599298
rect 157266 599144 177062 599298
rect 177230 599144 197670 599298
rect 197838 599144 217634 599298
rect 217802 599144 237598 599298
rect 237766 599144 258206 599298
rect 258374 599144 278170 599298
rect 278338 599144 298134 599298
rect 298302 599144 318742 599298
rect 318910 599144 338706 599298
rect 338874 599144 358670 599298
rect 358838 599144 379278 599298
rect 379446 599144 399242 599298
rect 399410 599144 419206 599298
rect 419374 599144 439814 599298
rect 439982 599144 459778 599298
rect 459946 599144 479742 599298
rect 479910 599144 499706 599298
rect 20 856 499816 599144
rect 130 734 19926 856
rect 20094 734 39890 856
rect 40058 734 59854 856
rect 60022 734 80462 856
rect 80630 734 100426 856
rect 100594 734 120390 856
rect 120558 734 140998 856
rect 141166 734 160962 856
rect 161130 734 180926 856
rect 181094 734 201534 856
rect 201702 734 221498 856
rect 221666 734 241462 856
rect 241630 734 262070 856
rect 262238 734 282034 856
rect 282202 734 301998 856
rect 302166 734 322606 856
rect 322774 734 342570 856
rect 342738 734 362534 856
rect 362702 734 383142 856
rect 383310 734 403106 856
rect 403274 734 423070 856
rect 423238 734 443678 856
rect 443846 734 463642 856
rect 463810 734 483606 856
rect 483774 734 499816 856
<< metal3 >>
rect 0 595688 800 595808
rect 499200 578688 500000 578808
rect 0 574608 800 574728
rect 499200 557608 500000 557728
rect 0 553528 800 553648
rect 499200 536528 500000 536648
rect 0 532448 800 532568
rect 499200 514768 500000 514888
rect 0 510688 800 510808
rect 499200 493688 500000 493808
rect 0 489608 800 489728
rect 499200 472608 500000 472728
rect 0 468528 800 468648
rect 499200 450848 500000 450968
rect 0 446768 800 446888
rect 499200 429768 500000 429888
rect 0 425688 800 425808
rect 499200 408688 500000 408808
rect 0 404608 800 404728
rect 499200 386928 500000 387048
rect 0 382848 800 382968
rect 499200 365848 500000 365968
rect 0 361768 800 361888
rect 499200 344768 500000 344888
rect 0 340688 800 340808
rect 499200 323008 500000 323128
rect 0 318928 800 319048
rect 499200 301928 500000 302048
rect 0 297848 800 297968
rect 499200 280848 500000 280968
rect 0 276768 800 276888
rect 499200 259088 500000 259208
rect 0 255008 800 255128
rect 499200 238008 500000 238128
rect 0 233928 800 234048
rect 499200 216928 500000 217048
rect 0 212848 800 212968
rect 499200 195168 500000 195288
rect 0 191088 800 191208
rect 499200 174088 500000 174208
rect 0 170008 800 170128
rect 499200 153008 500000 153128
rect 0 148928 800 149048
rect 499200 131248 500000 131368
rect 0 127168 800 127288
rect 499200 110168 500000 110288
rect 0 106088 800 106208
rect 499200 89088 500000 89208
rect 0 85008 800 85128
rect 499200 67328 500000 67448
rect 0 63248 800 63368
rect 499200 46248 500000 46368
rect 0 42168 800 42288
rect 499200 25168 500000 25288
rect 0 21088 800 21208
rect 499200 4088 500000 4208
<< obsm3 >>
rect 798 595888 499200 597345
rect 880 595608 499200 595888
rect 798 578888 499200 595608
rect 798 578608 499120 578888
rect 798 574808 499200 578608
rect 880 574528 499200 574808
rect 798 557808 499200 574528
rect 798 557528 499120 557808
rect 798 553728 499200 557528
rect 880 553448 499200 553728
rect 798 536728 499200 553448
rect 798 536448 499120 536728
rect 798 532648 499200 536448
rect 880 532368 499200 532648
rect 798 514968 499200 532368
rect 798 514688 499120 514968
rect 798 510888 499200 514688
rect 880 510608 499200 510888
rect 798 493888 499200 510608
rect 798 493608 499120 493888
rect 798 489808 499200 493608
rect 880 489528 499200 489808
rect 798 472808 499200 489528
rect 798 472528 499120 472808
rect 798 468728 499200 472528
rect 880 468448 499200 468728
rect 798 451048 499200 468448
rect 798 450768 499120 451048
rect 798 446968 499200 450768
rect 880 446688 499200 446968
rect 798 429968 499200 446688
rect 798 429688 499120 429968
rect 798 425888 499200 429688
rect 880 425608 499200 425888
rect 798 408888 499200 425608
rect 798 408608 499120 408888
rect 798 404808 499200 408608
rect 880 404528 499200 404808
rect 798 387128 499200 404528
rect 798 386848 499120 387128
rect 798 383048 499200 386848
rect 880 382768 499200 383048
rect 798 366048 499200 382768
rect 798 365768 499120 366048
rect 798 361968 499200 365768
rect 880 361688 499200 361968
rect 798 344968 499200 361688
rect 798 344688 499120 344968
rect 798 340888 499200 344688
rect 880 340608 499200 340888
rect 798 323208 499200 340608
rect 798 322928 499120 323208
rect 798 319128 499200 322928
rect 880 318848 499200 319128
rect 798 302128 499200 318848
rect 798 301848 499120 302128
rect 798 298048 499200 301848
rect 880 297768 499200 298048
rect 798 281048 499200 297768
rect 798 280768 499120 281048
rect 798 276968 499200 280768
rect 880 276688 499200 276968
rect 798 259288 499200 276688
rect 798 259008 499120 259288
rect 798 255208 499200 259008
rect 880 254928 499200 255208
rect 798 238208 499200 254928
rect 798 237928 499120 238208
rect 798 234128 499200 237928
rect 880 233848 499200 234128
rect 798 217128 499200 233848
rect 798 216848 499120 217128
rect 798 213048 499200 216848
rect 880 212768 499200 213048
rect 798 195368 499200 212768
rect 798 195088 499120 195368
rect 798 191288 499200 195088
rect 880 191008 499200 191288
rect 798 174288 499200 191008
rect 798 174008 499120 174288
rect 798 170208 499200 174008
rect 880 169928 499200 170208
rect 798 153208 499200 169928
rect 798 152928 499120 153208
rect 798 149128 499200 152928
rect 880 148848 499200 149128
rect 798 131448 499200 148848
rect 798 131168 499120 131448
rect 798 127368 499200 131168
rect 880 127088 499200 127368
rect 798 110368 499200 127088
rect 798 110088 499120 110368
rect 798 106288 499200 110088
rect 880 106008 499200 106288
rect 798 89288 499200 106008
rect 798 89008 499120 89288
rect 798 85208 499200 89008
rect 880 84928 499200 85208
rect 798 67528 499200 84928
rect 798 67248 499120 67528
rect 798 63448 499200 67248
rect 880 63168 499200 63448
rect 798 46448 499200 63168
rect 798 46168 499120 46448
rect 798 42368 499200 46168
rect 880 42088 499200 42368
rect 798 25368 499200 42088
rect 798 25088 499120 25368
rect 798 21288 499200 25088
rect 880 21008 499200 21288
rect 798 4288 499200 21008
rect 798 4008 499120 4288
rect 798 2143 499200 4008
<< metal4 >>
rect 4208 2128 4528 597360
rect 19568 2128 19888 597360
rect 34928 2128 35248 597360
rect 50288 2128 50608 597360
rect 65648 2128 65968 597360
rect 81008 2128 81328 597360
rect 96368 2128 96688 597360
rect 111728 2128 112048 597360
rect 127088 2128 127408 597360
rect 142448 2128 142768 597360
rect 157808 2128 158128 597360
rect 173168 2128 173488 597360
rect 188528 2128 188848 597360
rect 203888 2128 204208 597360
rect 219248 2128 219568 597360
rect 234608 2128 234928 597360
rect 249968 2128 250288 597360
rect 265328 2128 265648 597360
rect 280688 2128 281008 597360
rect 296048 2128 296368 597360
rect 311408 2128 311728 597360
rect 326768 2128 327088 597360
rect 342128 2128 342448 597360
rect 357488 2128 357808 597360
rect 372848 2128 373168 597360
rect 388208 2128 388528 597360
rect 403568 2128 403888 597360
rect 418928 2128 419248 597360
rect 434288 2128 434608 597360
rect 449648 2128 449968 597360
rect 465008 2128 465328 597360
rect 480368 2128 480688 597360
rect 495728 2128 496048 597360
<< obsm4 >>
rect 116347 2347 127008 597141
rect 127488 2347 142368 597141
rect 142848 2347 157728 597141
rect 158208 2347 173088 597141
rect 173568 2347 188448 597141
rect 188928 2347 203808 597141
rect 204288 2347 219168 597141
rect 219648 2347 234528 597141
rect 235008 2347 249888 597141
rect 250368 2347 265248 597141
rect 265728 2347 280608 597141
rect 281088 2347 295968 597141
rect 296448 2347 311328 597141
rect 311808 2347 326688 597141
rect 327168 2347 342048 597141
rect 342528 2347 357408 597141
rect 357888 2347 372768 597141
rect 373248 2347 373645 597141
<< labels >>
rlabel metal2 s 16118 599200 16174 600000 6 clk
port 1 nsew signal input
rlabel metal2 s 483662 0 483718 800 6 rst
port 2 nsew signal input
rlabel metal4 s 4208 2128 4528 597360 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 597360 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 597360 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 597360 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 597360 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 597360 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 597360 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 597360 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 597360 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 597360 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 597360 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 597360 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 597360 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 597360 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 597360 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 597360 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 597360 6 vccd1
port 3 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 597360 6 vssd1
port 4 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 597360 6 vssd1
port 4 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 597360 6 vssd1
port 4 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 597360 6 vssd1
port 4 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 597360 6 vssd1
port 4 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 597360 6 vssd1
port 4 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 597360 6 vssd1
port 4 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 597360 6 vssd1
port 4 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 597360 6 vssd1
port 4 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 597360 6 vssd1
port 4 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 597360 6 vssd1
port 4 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 597360 6 vssd1
port 4 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 597360 6 vssd1
port 4 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 597360 6 vssd1
port 4 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 597360 6 vssd1
port 4 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 597360 6 vssd1
port 4 nsew ground bidirectional
rlabel metal3 s 499200 493688 500000 493808 6 wbs_ack_o
port 5 nsew signal output
rlabel metal3 s 0 318928 800 319048 6 wbs_adr_i[0]
port 6 nsew signal input
rlabel metal3 s 0 361768 800 361888 6 wbs_adr_i[10]
port 7 nsew signal input
rlabel metal2 s 298190 599200 298246 600000 6 wbs_adr_i[11]
port 8 nsew signal input
rlabel metal2 s 358726 599200 358782 600000 6 wbs_adr_i[12]
port 9 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 wbs_adr_i[13]
port 10 nsew signal input
rlabel metal3 s 0 255008 800 255128 6 wbs_adr_i[14]
port 11 nsew signal input
rlabel metal3 s 499200 429768 500000 429888 6 wbs_adr_i[15]
port 12 nsew signal input
rlabel metal3 s 499200 344768 500000 344888 6 wbs_adr_i[16]
port 13 nsew signal input
rlabel metal3 s 499200 67328 500000 67448 6 wbs_adr_i[17]
port 14 nsew signal input
rlabel metal3 s 0 425688 800 425808 6 wbs_adr_i[18]
port 15 nsew signal input
rlabel metal2 s 342626 0 342682 800 6 wbs_adr_i[19]
port 16 nsew signal input
rlabel metal2 s 463698 0 463754 800 6 wbs_adr_i[1]
port 17 nsew signal input
rlabel metal3 s 499200 174088 500000 174208 6 wbs_adr_i[20]
port 18 nsew signal input
rlabel metal2 s 237654 599200 237710 600000 6 wbs_adr_i[21]
port 19 nsew signal input
rlabel metal3 s 0 468528 800 468648 6 wbs_adr_i[22]
port 20 nsew signal input
rlabel metal2 s 116582 599200 116638 600000 6 wbs_adr_i[23]
port 21 nsew signal input
rlabel metal3 s 499200 557608 500000 557728 6 wbs_adr_i[24]
port 22 nsew signal input
rlabel metal2 s 278226 599200 278282 600000 6 wbs_adr_i[25]
port 23 nsew signal input
rlabel metal3 s 499200 153008 500000 153128 6 wbs_adr_i[26]
port 24 nsew signal input
rlabel metal3 s 0 297848 800 297968 6 wbs_adr_i[27]
port 25 nsew signal input
rlabel metal2 s 221554 0 221610 800 6 wbs_adr_i[28]
port 26 nsew signal input
rlabel metal3 s 0 191088 800 191208 6 wbs_adr_i[29]
port 27 nsew signal input
rlabel metal3 s 499200 131248 500000 131368 6 wbs_adr_i[2]
port 28 nsew signal input
rlabel metal2 s 338762 599200 338818 600000 6 wbs_adr_i[30]
port 29 nsew signal input
rlabel metal3 s 0 382848 800 382968 6 wbs_adr_i[31]
port 30 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 wbs_adr_i[3]
port 31 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 wbs_adr_i[4]
port 32 nsew signal input
rlabel metal2 s 459834 599200 459890 600000 6 wbs_adr_i[5]
port 33 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 wbs_adr_i[6]
port 34 nsew signal input
rlabel metal3 s 0 106088 800 106208 6 wbs_adr_i[7]
port 35 nsew signal input
rlabel metal2 s 499762 599200 499818 600000 6 wbs_adr_i[8]
port 36 nsew signal input
rlabel metal2 s 399298 599200 399354 600000 6 wbs_adr_i[9]
port 37 nsew signal input
rlabel metal3 s 499200 514768 500000 514888 6 wbs_cyc_i
port 38 nsew signal input
rlabel metal3 s 499200 578688 500000 578808 6 wbs_dat_i[0]
port 39 nsew signal input
rlabel metal3 s 499200 280848 500000 280968 6 wbs_dat_i[10]
port 40 nsew signal input
rlabel metal3 s 499200 238008 500000 238128 6 wbs_dat_i[11]
port 41 nsew signal input
rlabel metal2 s 137190 599200 137246 600000 6 wbs_dat_i[12]
port 42 nsew signal input
rlabel metal2 s 157154 599200 157210 600000 6 wbs_dat_i[13]
port 43 nsew signal input
rlabel metal3 s 499200 472608 500000 472728 6 wbs_dat_i[14]
port 44 nsew signal input
rlabel metal2 s 217690 599200 217746 600000 6 wbs_dat_i[15]
port 45 nsew signal input
rlabel metal2 s 141054 0 141110 800 6 wbs_dat_i[16]
port 46 nsew signal input
rlabel metal2 s 177118 599200 177174 600000 6 wbs_dat_i[17]
port 47 nsew signal input
rlabel metal3 s 499200 46248 500000 46368 6 wbs_dat_i[18]
port 48 nsew signal input
rlabel metal2 s 258262 599200 258318 600000 6 wbs_dat_i[19]
port 49 nsew signal input
rlabel metal3 s 0 404608 800 404728 6 wbs_dat_i[1]
port 50 nsew signal input
rlabel metal2 s 96618 599200 96674 600000 6 wbs_dat_i[20]
port 51 nsew signal input
rlabel metal3 s 499200 89088 500000 89208 6 wbs_dat_i[21]
port 52 nsew signal input
rlabel metal3 s 499200 536528 500000 536648 6 wbs_dat_i[22]
port 53 nsew signal input
rlabel metal2 s 419262 599200 419318 600000 6 wbs_dat_i[23]
port 54 nsew signal input
rlabel metal2 s 403162 0 403218 800 6 wbs_dat_i[24]
port 55 nsew signal input
rlabel metal2 s 201590 0 201646 800 6 wbs_dat_i[25]
port 56 nsew signal input
rlabel metal3 s 499200 195168 500000 195288 6 wbs_dat_i[26]
port 57 nsew signal input
rlabel metal3 s 0 212848 800 212968 6 wbs_dat_i[27]
port 58 nsew signal input
rlabel metal3 s 0 276768 800 276888 6 wbs_dat_i[28]
port 59 nsew signal input
rlabel metal3 s 499200 25168 500000 25288 6 wbs_dat_i[29]
port 60 nsew signal input
rlabel metal2 s 56046 599200 56102 600000 6 wbs_dat_i[2]
port 61 nsew signal input
rlabel metal2 s 423126 0 423182 800 6 wbs_dat_i[30]
port 62 nsew signal input
rlabel metal3 s 0 510688 800 510808 6 wbs_dat_i[31]
port 63 nsew signal input
rlabel metal3 s 0 85008 800 85128 6 wbs_dat_i[3]
port 64 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 wbs_dat_i[4]
port 65 nsew signal input
rlabel metal2 s 161018 0 161074 800 6 wbs_dat_i[5]
port 66 nsew signal input
rlabel metal3 s 499200 4088 500000 4208 6 wbs_dat_i[6]
port 67 nsew signal input
rlabel metal3 s 499200 323008 500000 323128 6 wbs_dat_i[7]
port 68 nsew signal input
rlabel metal3 s 499200 216928 500000 217048 6 wbs_dat_i[8]
port 69 nsew signal input
rlabel metal2 s 383198 0 383254 800 6 wbs_dat_i[9]
port 70 nsew signal input
rlabel metal3 s 0 446768 800 446888 6 wbs_dat_o[0]
port 71 nsew signal output
rlabel metal3 s 0 340688 800 340808 6 wbs_dat_o[10]
port 72 nsew signal output
rlabel metal3 s 0 127168 800 127288 6 wbs_dat_o[11]
port 73 nsew signal output
rlabel metal3 s 499200 259088 500000 259208 6 wbs_dat_o[12]
port 74 nsew signal output
rlabel metal3 s 499200 408688 500000 408808 6 wbs_dat_o[13]
port 75 nsew signal output
rlabel metal2 s 443734 0 443790 800 6 wbs_dat_o[14]
port 76 nsew signal output
rlabel metal3 s 499200 450848 500000 450968 6 wbs_dat_o[15]
port 77 nsew signal output
rlabel metal2 s 262126 0 262182 800 6 wbs_dat_o[16]
port 78 nsew signal output
rlabel metal3 s 0 553528 800 553648 6 wbs_dat_o[17]
port 79 nsew signal output
rlabel metal3 s 0 233928 800 234048 6 wbs_dat_o[18]
port 80 nsew signal output
rlabel metal2 s 18 0 74 800 6 wbs_dat_o[19]
port 81 nsew signal output
rlabel metal2 s 322662 0 322718 800 6 wbs_dat_o[1]
port 82 nsew signal output
rlabel metal2 s 36082 599200 36138 600000 6 wbs_dat_o[20]
port 83 nsew signal output
rlabel metal2 s 197726 599200 197782 600000 6 wbs_dat_o[21]
port 84 nsew signal output
rlabel metal3 s 0 63248 800 63368 6 wbs_dat_o[22]
port 85 nsew signal output
rlabel metal3 s 0 532448 800 532568 6 wbs_dat_o[23]
port 86 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 wbs_dat_o[24]
port 87 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_o[25]
port 88 nsew signal output
rlabel metal2 s 439870 599200 439926 600000 6 wbs_dat_o[26]
port 89 nsew signal output
rlabel metal2 s 318798 599200 318854 600000 6 wbs_dat_o[27]
port 90 nsew signal output
rlabel metal2 s 241518 0 241574 800 6 wbs_dat_o[28]
port 91 nsew signal output
rlabel metal2 s 479798 599200 479854 600000 6 wbs_dat_o[29]
port 92 nsew signal output
rlabel metal3 s 499200 110168 500000 110288 6 wbs_dat_o[2]
port 93 nsew signal output
rlabel metal3 s 0 574608 800 574728 6 wbs_dat_o[30]
port 94 nsew signal output
rlabel metal3 s 499200 365848 500000 365968 6 wbs_dat_o[31]
port 95 nsew signal output
rlabel metal2 s 100482 0 100538 800 6 wbs_dat_o[3]
port 96 nsew signal output
rlabel metal2 s 180982 0 181038 800 6 wbs_dat_o[4]
port 97 nsew signal output
rlabel metal2 s 282090 0 282146 800 6 wbs_dat_o[5]
port 98 nsew signal output
rlabel metal3 s 499200 386928 500000 387048 6 wbs_dat_o[6]
port 99 nsew signal output
rlabel metal2 s 302054 0 302110 800 6 wbs_dat_o[7]
port 100 nsew signal output
rlabel metal3 s 0 148928 800 149048 6 wbs_dat_o[8]
port 101 nsew signal output
rlabel metal2 s 379334 599200 379390 600000 6 wbs_dat_o[9]
port 102 nsew signal output
rlabel metal3 s 0 595688 800 595808 6 wbs_sel_i[0]
port 103 nsew signal input
rlabel metal2 s 76654 599200 76710 600000 6 wbs_sel_i[1]
port 104 nsew signal input
rlabel metal2 s 362590 0 362646 800 6 wbs_sel_i[2]
port 105 nsew signal input
rlabel metal3 s 0 170008 800 170128 6 wbs_sel_i[3]
port 106 nsew signal input
rlabel metal3 s 0 489608 800 489728 6 wbs_stb_i
port 107 nsew signal input
rlabel metal3 s 499200 301928 500000 302048 6 wbs_we_i
port 108 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 500000 600000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 274525888
string GDS_FILE /home/edabk/efabless/caravel_user_project/openlane/neuron_core/runs/23_11_06_07_26/results/signoff/neuron_core.magic.gds
string GDS_START 1565098
<< end >>

