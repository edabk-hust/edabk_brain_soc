version https://git-lfs.github.com/spec/v1
oid sha256:5e0c79900648c1b3513bccb333bb8f73ea3e3130a7fd0d3721ee1de68ad07c2f
size 163323
