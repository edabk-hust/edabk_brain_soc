version https://git-lfs.github.com/spec/v1
oid sha256:6adbc7cca35d4c1a802eb07682d4d5cfbb3d8f540b7585e697c999af414f6159
size 59743791
